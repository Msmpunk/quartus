library ieee;
use ieee.std_logic_1164.all;
entity xorproject is
port(
a,b: in std_logic;

c:out std_logic);
end;

architecture arqxorproject of xorproject is
begin
c<= a xor b;
end;